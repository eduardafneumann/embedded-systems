// SEProjetoFinalSingle.v

// Generated using ACDS version 21.1 850

`timescale 1 ps / 1 ps
module SEProjetoFinalSingle (
		input  wire  clk_clk  // clk.clk
	);

	wire         cpu0_debug_reset_request_reset;                        // CPU0:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] cpu0_data_master_readdata;                             // mm_interconnect_0:CPU0_data_master_readdata -> CPU0:d_readdata
	wire         cpu0_data_master_waitrequest;                          // mm_interconnect_0:CPU0_data_master_waitrequest -> CPU0:d_waitrequest
	wire         cpu0_data_master_debugaccess;                          // CPU0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU0_data_master_debugaccess
	wire  [19:0] cpu0_data_master_address;                              // CPU0:d_address -> mm_interconnect_0:CPU0_data_master_address
	wire   [3:0] cpu0_data_master_byteenable;                           // CPU0:d_byteenable -> mm_interconnect_0:CPU0_data_master_byteenable
	wire         cpu0_data_master_read;                                 // CPU0:d_read -> mm_interconnect_0:CPU0_data_master_read
	wire         cpu0_data_master_readdatavalid;                        // mm_interconnect_0:CPU0_data_master_readdatavalid -> CPU0:d_readdatavalid
	wire         cpu0_data_master_write;                                // CPU0:d_write -> mm_interconnect_0:CPU0_data_master_write
	wire  [31:0] cpu0_data_master_writedata;                            // CPU0:d_writedata -> mm_interconnect_0:CPU0_data_master_writedata
	wire  [31:0] cpu0_instruction_master_readdata;                      // mm_interconnect_0:CPU0_instruction_master_readdata -> CPU0:i_readdata
	wire         cpu0_instruction_master_waitrequest;                   // mm_interconnect_0:CPU0_instruction_master_waitrequest -> CPU0:i_waitrequest
	wire  [19:0] cpu0_instruction_master_address;                       // CPU0:i_address -> mm_interconnect_0:CPU0_instruction_master_address
	wire         cpu0_instruction_master_read;                          // CPU0:i_read -> mm_interconnect_0:CPU0_instruction_master_read
	wire         cpu0_instruction_master_readdatavalid;                 // mm_interconnect_0:CPU0_instruction_master_readdatavalid -> CPU0:i_readdatavalid
	wire         mm_interconnect_0_uart0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:UART0_avalon_jtag_slave_chipselect -> UART0:av_chipselect
	wire  [31:0] mm_interconnect_0_uart0_avalon_jtag_slave_readdata;    // UART0:av_readdata -> mm_interconnect_0:UART0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_uart0_avalon_jtag_slave_waitrequest; // UART0:av_waitrequest -> mm_interconnect_0:UART0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_uart0_avalon_jtag_slave_address;     // mm_interconnect_0:UART0_avalon_jtag_slave_address -> UART0:av_address
	wire         mm_interconnect_0_uart0_avalon_jtag_slave_read;        // mm_interconnect_0:UART0_avalon_jtag_slave_read -> UART0:av_read_n
	wire         mm_interconnect_0_uart0_avalon_jtag_slave_write;       // mm_interconnect_0:UART0_avalon_jtag_slave_write -> UART0:av_write_n
	wire  [31:0] mm_interconnect_0_uart0_avalon_jtag_slave_writedata;   // mm_interconnect_0:UART0_avalon_jtag_slave_writedata -> UART0:av_writedata
	wire  [31:0] mm_interconnect_0_cpu0_debug_mem_slave_readdata;       // CPU0:debug_mem_slave_readdata -> mm_interconnect_0:CPU0_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu0_debug_mem_slave_waitrequest;    // CPU0:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu0_debug_mem_slave_debugaccess;    // mm_interconnect_0:CPU0_debug_mem_slave_debugaccess -> CPU0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu0_debug_mem_slave_address;        // mm_interconnect_0:CPU0_debug_mem_slave_address -> CPU0:debug_mem_slave_address
	wire         mm_interconnect_0_cpu0_debug_mem_slave_read;           // mm_interconnect_0:CPU0_debug_mem_slave_read -> CPU0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu0_debug_mem_slave_byteenable;     // mm_interconnect_0:CPU0_debug_mem_slave_byteenable -> CPU0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu0_debug_mem_slave_write;          // mm_interconnect_0:CPU0_debug_mem_slave_write -> CPU0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu0_debug_mem_slave_writedata;      // mm_interconnect_0:CPU0_debug_mem_slave_writedata -> CPU0:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                 // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:chipselect
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                   // SDRAM:readdata -> mm_interconnect_0:SDRAM_s1_readdata
	wire  [15:0] mm_interconnect_0_sdram_s1_address;                    // mm_interconnect_0:SDRAM_s1_address -> SDRAM:address
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                 // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:byteenable
	wire         mm_interconnect_0_sdram_s1_write;                      // mm_interconnect_0:SDRAM_s1_write -> SDRAM:write
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                  // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:writedata
	wire         mm_interconnect_0_sdram_s1_clken;                      // mm_interconnect_0:SDRAM_s1_clken -> SDRAM:clken
	wire         irq_mapper_receiver0_irq;                              // UART0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu0_irq_irq;                                          // irq_mapper:sender_irq -> CPU0:irq
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [CPU0:reset_n, SDRAM:reset, UART0:rst_n, irq_mapper:reset, mm_interconnect_0:CPU0_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                    // rst_controller:reset_req -> [CPU0:reset_req, SDRAM:reset_req, rst_translator:reset_req_in]

	SEProjetoFinalSingle_CPU0 cpu0 (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (cpu0_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu0_data_master_read),                              //                          .read
		.d_readdata                          (cpu0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu0_data_master_write),                             //                          .write
		.d_writedata                         (cpu0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu0_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	SEProjetoFinalSingle_SDRAM sdram (
		.clk        (clk_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_sdram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sdram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sdram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sdram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sdram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sdram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sdram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze     (1'b0)                                   // (terminated)
	);

	SEProjetoFinalSingle_UART0 uart0 (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_uart0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_uart0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_uart0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_uart0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_uart0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_uart0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_uart0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                               //               irq.irq
	);

	SEProjetoFinalSingle_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                          (clk_clk),                                               //                        clk_0_clk.clk
		.CPU0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // CPU0_reset_reset_bridge_in_reset.reset
		.CPU0_data_master_address               (cpu0_data_master_address),                              //                 CPU0_data_master.address
		.CPU0_data_master_waitrequest           (cpu0_data_master_waitrequest),                          //                                 .waitrequest
		.CPU0_data_master_byteenable            (cpu0_data_master_byteenable),                           //                                 .byteenable
		.CPU0_data_master_read                  (cpu0_data_master_read),                                 //                                 .read
		.CPU0_data_master_readdata              (cpu0_data_master_readdata),                             //                                 .readdata
		.CPU0_data_master_readdatavalid         (cpu0_data_master_readdatavalid),                        //                                 .readdatavalid
		.CPU0_data_master_write                 (cpu0_data_master_write),                                //                                 .write
		.CPU0_data_master_writedata             (cpu0_data_master_writedata),                            //                                 .writedata
		.CPU0_data_master_debugaccess           (cpu0_data_master_debugaccess),                          //                                 .debugaccess
		.CPU0_instruction_master_address        (cpu0_instruction_master_address),                       //          CPU0_instruction_master.address
		.CPU0_instruction_master_waitrequest    (cpu0_instruction_master_waitrequest),                   //                                 .waitrequest
		.CPU0_instruction_master_read           (cpu0_instruction_master_read),                          //                                 .read
		.CPU0_instruction_master_readdata       (cpu0_instruction_master_readdata),                      //                                 .readdata
		.CPU0_instruction_master_readdatavalid  (cpu0_instruction_master_readdatavalid),                 //                                 .readdatavalid
		.CPU0_debug_mem_slave_address           (mm_interconnect_0_cpu0_debug_mem_slave_address),        //             CPU0_debug_mem_slave.address
		.CPU0_debug_mem_slave_write             (mm_interconnect_0_cpu0_debug_mem_slave_write),          //                                 .write
		.CPU0_debug_mem_slave_read              (mm_interconnect_0_cpu0_debug_mem_slave_read),           //                                 .read
		.CPU0_debug_mem_slave_readdata          (mm_interconnect_0_cpu0_debug_mem_slave_readdata),       //                                 .readdata
		.CPU0_debug_mem_slave_writedata         (mm_interconnect_0_cpu0_debug_mem_slave_writedata),      //                                 .writedata
		.CPU0_debug_mem_slave_byteenable        (mm_interconnect_0_cpu0_debug_mem_slave_byteenable),     //                                 .byteenable
		.CPU0_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu0_debug_mem_slave_waitrequest),    //                                 .waitrequest
		.CPU0_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu0_debug_mem_slave_debugaccess),    //                                 .debugaccess
		.SDRAM_s1_address                       (mm_interconnect_0_sdram_s1_address),                    //                         SDRAM_s1.address
		.SDRAM_s1_write                         (mm_interconnect_0_sdram_s1_write),                      //                                 .write
		.SDRAM_s1_readdata                      (mm_interconnect_0_sdram_s1_readdata),                   //                                 .readdata
		.SDRAM_s1_writedata                     (mm_interconnect_0_sdram_s1_writedata),                  //                                 .writedata
		.SDRAM_s1_byteenable                    (mm_interconnect_0_sdram_s1_byteenable),                 //                                 .byteenable
		.SDRAM_s1_chipselect                    (mm_interconnect_0_sdram_s1_chipselect),                 //                                 .chipselect
		.SDRAM_s1_clken                         (mm_interconnect_0_sdram_s1_clken),                      //                                 .clken
		.UART0_avalon_jtag_slave_address        (mm_interconnect_0_uart0_avalon_jtag_slave_address),     //          UART0_avalon_jtag_slave.address
		.UART0_avalon_jtag_slave_write          (mm_interconnect_0_uart0_avalon_jtag_slave_write),       //                                 .write
		.UART0_avalon_jtag_slave_read           (mm_interconnect_0_uart0_avalon_jtag_slave_read),        //                                 .read
		.UART0_avalon_jtag_slave_readdata       (mm_interconnect_0_uart0_avalon_jtag_slave_readdata),    //                                 .readdata
		.UART0_avalon_jtag_slave_writedata      (mm_interconnect_0_uart0_avalon_jtag_slave_writedata),   //                                 .writedata
		.UART0_avalon_jtag_slave_waitrequest    (mm_interconnect_0_uart0_avalon_jtag_slave_waitrequest), //                                 .waitrequest
		.UART0_avalon_jtag_slave_chipselect     (mm_interconnect_0_uart0_avalon_jtag_slave_chipselect)   //                                 .chipselect
	);

	SEProjetoFinalSingle_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu0_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (cpu0_debug_reset_request_reset),     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
