
module SEProjetoFinal (
	clk_clk);	

	input		clk_clk;
endmodule
