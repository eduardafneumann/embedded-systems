// SEProjetoFinal.v

// Generated using ACDS version 21.1 850

`timescale 1 ps / 1 ps
module SEProjetoFinal (
		input  wire  clk_clk  // clk.clk
	);

	wire         cpu0_debug_reset_request_reset;                     // CPU0:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] cpu0_data_master_readdata;                          // mm_interconnect_0:CPU0_data_master_readdata -> CPU0:d_readdata
	wire         cpu0_data_master_waitrequest;                       // mm_interconnect_0:CPU0_data_master_waitrequest -> CPU0:d_waitrequest
	wire         cpu0_data_master_debugaccess;                       // CPU0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU0_data_master_debugaccess
	wire  [18:0] cpu0_data_master_address;                           // CPU0:d_address -> mm_interconnect_0:CPU0_data_master_address
	wire   [3:0] cpu0_data_master_byteenable;                        // CPU0:d_byteenable -> mm_interconnect_0:CPU0_data_master_byteenable
	wire         cpu0_data_master_read;                              // CPU0:d_read -> mm_interconnect_0:CPU0_data_master_read
	wire         cpu0_data_master_readdatavalid;                     // mm_interconnect_0:CPU0_data_master_readdatavalid -> CPU0:d_readdatavalid
	wire         cpu0_data_master_write;                             // CPU0:d_write -> mm_interconnect_0:CPU0_data_master_write
	wire  [31:0] cpu0_data_master_writedata;                         // CPU0:d_writedata -> mm_interconnect_0:CPU0_data_master_writedata
	wire  [31:0] cpu0_instruction_master_readdata;                   // mm_interconnect_0:CPU0_instruction_master_readdata -> CPU0:i_readdata
	wire         cpu0_instruction_master_waitrequest;                // mm_interconnect_0:CPU0_instruction_master_waitrequest -> CPU0:i_waitrequest
	wire  [18:0] cpu0_instruction_master_address;                    // CPU0:i_address -> mm_interconnect_0:CPU0_instruction_master_address
	wire         cpu0_instruction_master_read;                       // CPU0:i_read -> mm_interconnect_0:CPU0_instruction_master_read
	wire         cpu0_instruction_master_readdatavalid;              // mm_interconnect_0:CPU0_instruction_master_readdatavalid -> CPU0:i_readdatavalid
	wire  [31:0] cpu1_data_master_readdata;                          // mm_interconnect_0:CPU1_data_master_readdata -> CPU1:d_readdata
	wire         cpu1_data_master_waitrequest;                       // mm_interconnect_0:CPU1_data_master_waitrequest -> CPU1:d_waitrequest
	wire         cpu1_data_master_debugaccess;                       // CPU1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU1_data_master_debugaccess
	wire  [18:0] cpu1_data_master_address;                           // CPU1:d_address -> mm_interconnect_0:CPU1_data_master_address
	wire   [3:0] cpu1_data_master_byteenable;                        // CPU1:d_byteenable -> mm_interconnect_0:CPU1_data_master_byteenable
	wire         cpu1_data_master_read;                              // CPU1:d_read -> mm_interconnect_0:CPU1_data_master_read
	wire         cpu1_data_master_readdatavalid;                     // mm_interconnect_0:CPU1_data_master_readdatavalid -> CPU1:d_readdatavalid
	wire         cpu1_data_master_write;                             // CPU1:d_write -> mm_interconnect_0:CPU1_data_master_write
	wire  [31:0] cpu1_data_master_writedata;                         // CPU1:d_writedata -> mm_interconnect_0:CPU1_data_master_writedata
	wire  [31:0] cpu2_data_master_readdata;                          // mm_interconnect_0:CPU2_data_master_readdata -> CPU2:d_readdata
	wire         cpu2_data_master_waitrequest;                       // mm_interconnect_0:CPU2_data_master_waitrequest -> CPU2:d_waitrequest
	wire         cpu2_data_master_debugaccess;                       // CPU2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU2_data_master_debugaccess
	wire  [18:0] cpu2_data_master_address;                           // CPU2:d_address -> mm_interconnect_0:CPU2_data_master_address
	wire   [3:0] cpu2_data_master_byteenable;                        // CPU2:d_byteenable -> mm_interconnect_0:CPU2_data_master_byteenable
	wire         cpu2_data_master_read;                              // CPU2:d_read -> mm_interconnect_0:CPU2_data_master_read
	wire         cpu2_data_master_readdatavalid;                     // mm_interconnect_0:CPU2_data_master_readdatavalid -> CPU2:d_readdatavalid
	wire         cpu2_data_master_write;                             // CPU2:d_write -> mm_interconnect_0:CPU2_data_master_write
	wire  [31:0] cpu2_data_master_writedata;                         // CPU2:d_writedata -> mm_interconnect_0:CPU2_data_master_writedata
	wire  [31:0] cpu3_data_master_readdata;                          // mm_interconnect_0:CPU3_data_master_readdata -> CPU3:d_readdata
	wire         cpu3_data_master_waitrequest;                       // mm_interconnect_0:CPU3_data_master_waitrequest -> CPU3:d_waitrequest
	wire         cpu3_data_master_debugaccess;                       // CPU3:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU3_data_master_debugaccess
	wire  [18:0] cpu3_data_master_address;                           // CPU3:d_address -> mm_interconnect_0:CPU3_data_master_address
	wire   [3:0] cpu3_data_master_byteenable;                        // CPU3:d_byteenable -> mm_interconnect_0:CPU3_data_master_byteenable
	wire         cpu3_data_master_read;                              // CPU3:d_read -> mm_interconnect_0:CPU3_data_master_read
	wire         cpu3_data_master_readdatavalid;                     // mm_interconnect_0:CPU3_data_master_readdatavalid -> CPU3:d_readdatavalid
	wire         cpu3_data_master_write;                             // CPU3:d_write -> mm_interconnect_0:CPU3_data_master_write
	wire  [31:0] cpu3_data_master_writedata;                         // CPU3:d_writedata -> mm_interconnect_0:CPU3_data_master_writedata
	wire  [31:0] cpu1_instruction_master_readdata;                   // mm_interconnect_0:CPU1_instruction_master_readdata -> CPU1:i_readdata
	wire         cpu1_instruction_master_waitrequest;                // mm_interconnect_0:CPU1_instruction_master_waitrequest -> CPU1:i_waitrequest
	wire  [18:0] cpu1_instruction_master_address;                    // CPU1:i_address -> mm_interconnect_0:CPU1_instruction_master_address
	wire         cpu1_instruction_master_read;                       // CPU1:i_read -> mm_interconnect_0:CPU1_instruction_master_read
	wire         cpu1_instruction_master_readdatavalid;              // mm_interconnect_0:CPU1_instruction_master_readdatavalid -> CPU1:i_readdatavalid
	wire  [31:0] cpu2_instruction_master_readdata;                   // mm_interconnect_0:CPU2_instruction_master_readdata -> CPU2:i_readdata
	wire         cpu2_instruction_master_waitrequest;                // mm_interconnect_0:CPU2_instruction_master_waitrequest -> CPU2:i_waitrequest
	wire  [18:0] cpu2_instruction_master_address;                    // CPU2:i_address -> mm_interconnect_0:CPU2_instruction_master_address
	wire         cpu2_instruction_master_read;                       // CPU2:i_read -> mm_interconnect_0:CPU2_instruction_master_read
	wire         cpu2_instruction_master_readdatavalid;              // mm_interconnect_0:CPU2_instruction_master_readdatavalid -> CPU2:i_readdatavalid
	wire  [31:0] cpu3_instruction_master_readdata;                   // mm_interconnect_0:CPU3_instruction_master_readdata -> CPU3:i_readdata
	wire         cpu3_instruction_master_waitrequest;                // mm_interconnect_0:CPU3_instruction_master_waitrequest -> CPU3:i_waitrequest
	wire  [18:0] cpu3_instruction_master_address;                    // CPU3:i_address -> mm_interconnect_0:CPU3_instruction_master_address
	wire         cpu3_instruction_master_read;                       // CPU3:i_read -> mm_interconnect_0:CPU3_instruction_master_read
	wire         cpu3_instruction_master_readdatavalid;              // mm_interconnect_0:CPU3_instruction_master_readdatavalid -> CPU3:i_readdatavalid
	wire  [31:0] mm_interconnect_0_cpu0_debug_mem_slave_readdata;    // CPU0:debug_mem_slave_readdata -> mm_interconnect_0:CPU0_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu0_debug_mem_slave_waitrequest; // CPU0:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu0_debug_mem_slave_debugaccess; // mm_interconnect_0:CPU0_debug_mem_slave_debugaccess -> CPU0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu0_debug_mem_slave_address;     // mm_interconnect_0:CPU0_debug_mem_slave_address -> CPU0:debug_mem_slave_address
	wire         mm_interconnect_0_cpu0_debug_mem_slave_read;        // mm_interconnect_0:CPU0_debug_mem_slave_read -> CPU0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu0_debug_mem_slave_byteenable;  // mm_interconnect_0:CPU0_debug_mem_slave_byteenable -> CPU0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu0_debug_mem_slave_write;       // mm_interconnect_0:CPU0_debug_mem_slave_write -> CPU0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu0_debug_mem_slave_writedata;   // mm_interconnect_0:CPU0_debug_mem_slave_writedata -> CPU0:debug_mem_slave_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;               // mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                 // SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	wire  [15:0] mm_interconnect_0_sram_s1_address;                  // mm_interconnect_0:SRAM_s1_address -> SRAM:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;               // mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_s1_write;                    // mm_interconnect_0:SRAM_s1_write -> SRAM:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                // mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	wire         mm_interconnect_0_sram_s1_clken;                    // mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	wire  [31:0] mm_interconnect_0_cpu3_debug_mem_slave_readdata;    // CPU3:debug_mem_slave_readdata -> mm_interconnect_0:CPU3_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu3_debug_mem_slave_waitrequest; // CPU3:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU3_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu3_debug_mem_slave_debugaccess; // mm_interconnect_0:CPU3_debug_mem_slave_debugaccess -> CPU3:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu3_debug_mem_slave_address;     // mm_interconnect_0:CPU3_debug_mem_slave_address -> CPU3:debug_mem_slave_address
	wire         mm_interconnect_0_cpu3_debug_mem_slave_read;        // mm_interconnect_0:CPU3_debug_mem_slave_read -> CPU3:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu3_debug_mem_slave_byteenable;  // mm_interconnect_0:CPU3_debug_mem_slave_byteenable -> CPU3:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu3_debug_mem_slave_write;       // mm_interconnect_0:CPU3_debug_mem_slave_write -> CPU3:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu3_debug_mem_slave_writedata;   // mm_interconnect_0:CPU3_debug_mem_slave_writedata -> CPU3:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_cpu2_debug_mem_slave_readdata;    // CPU2:debug_mem_slave_readdata -> mm_interconnect_0:CPU2_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu2_debug_mem_slave_waitrequest; // CPU2:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu2_debug_mem_slave_debugaccess; // mm_interconnect_0:CPU2_debug_mem_slave_debugaccess -> CPU2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu2_debug_mem_slave_address;     // mm_interconnect_0:CPU2_debug_mem_slave_address -> CPU2:debug_mem_slave_address
	wire         mm_interconnect_0_cpu2_debug_mem_slave_read;        // mm_interconnect_0:CPU2_debug_mem_slave_read -> CPU2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu2_debug_mem_slave_byteenable;  // mm_interconnect_0:CPU2_debug_mem_slave_byteenable -> CPU2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu2_debug_mem_slave_write;       // mm_interconnect_0:CPU2_debug_mem_slave_write -> CPU2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu2_debug_mem_slave_writedata;   // mm_interconnect_0:CPU2_debug_mem_slave_writedata -> CPU2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_cpu1_debug_mem_slave_readdata;    // CPU1:debug_mem_slave_readdata -> mm_interconnect_0:CPU1_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu1_debug_mem_slave_waitrequest; // CPU1:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU1_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu1_debug_mem_slave_debugaccess; // mm_interconnect_0:CPU1_debug_mem_slave_debugaccess -> CPU1:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu1_debug_mem_slave_address;     // mm_interconnect_0:CPU1_debug_mem_slave_address -> CPU1:debug_mem_slave_address
	wire         mm_interconnect_0_cpu1_debug_mem_slave_read;        // mm_interconnect_0:CPU1_debug_mem_slave_read -> CPU1:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu1_debug_mem_slave_byteenable;  // mm_interconnect_0:CPU1_debug_mem_slave_byteenable -> CPU1:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu1_debug_mem_slave_write;       // mm_interconnect_0:CPU1_debug_mem_slave_write -> CPU1:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu1_debug_mem_slave_writedata;   // mm_interconnect_0:CPU1_debug_mem_slave_writedata -> CPU1:debug_mem_slave_writedata
	wire         irq_mapper_receiver0_irq;                           // DEBUG:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu0_irq_irq;                                       // irq_mapper:sender_irq -> CPU0:irq
	wire  [31:0] cpu1_irq_irq;                                       // irq_mapper_001:sender_irq -> CPU1:irq
	wire  [31:0] cpu2_irq_irq;                                       // irq_mapper_002:sender_irq -> CPU2:irq
	wire  [31:0] cpu3_irq_irq;                                       // irq_mapper_003:sender_irq -> CPU3:irq
	wire         rst_controller_reset_out_reset;                     // rst_controller:reset_out -> [CPU0:reset_n, CPU1:reset_n, CPU2:reset_n, CPU3:reset_n, DEBUG:rst_n, SRAM:reset, irq_mapper:reset, irq_mapper_001:reset, irq_mapper_002:reset, irq_mapper_003:reset, mm_interconnect_0:CPU0_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                 // rst_controller:reset_req -> [CPU0:reset_req, CPU1:reset_req, CPU2:reset_req, CPU3:reset_req, SRAM:reset_req, rst_translator:reset_req_in]

	SEProjetoFinal_CPU0 cpu0 (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (cpu0_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu0_data_master_read),                              //                          .read
		.d_readdata                          (cpu0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu0_data_master_write),                             //                          .write
		.d_writedata                         (cpu0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu0_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	SEProjetoFinal_CPU1 cpu1 (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (cpu1_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu1_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu1_data_master_read),                              //                          .read
		.d_readdata                          (cpu1_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu1_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu1_data_master_write),                             //                          .write
		.d_writedata                         (cpu1_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu1_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu1_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu1_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu1_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu1_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu1_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu1_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu1_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                   //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu1_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu1_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu1_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu1_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu1_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu1_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu1_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu1_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	SEProjetoFinal_CPU2 cpu2 (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (cpu2_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu2_data_master_read),                              //                          .read
		.d_readdata                          (cpu2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu2_data_master_write),                             //                          .write
		.d_writedata                         (cpu2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu2_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                   //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	SEProjetoFinal_CPU3 cpu3 (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (cpu3_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu3_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu3_data_master_read),                              //                          .read
		.d_readdata                          (cpu3_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu3_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu3_data_master_write),                             //                          .write
		.d_writedata                         (cpu3_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu3_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu3_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu3_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu3_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu3_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu3_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu3_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu3_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                   //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu3_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu3_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu3_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu3_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu3_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu3_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu3_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu3_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	SEProjetoFinal_DEBUG debug (
		.clk            (clk_clk),                         //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset), //             reset.reset_n
		.av_chipselect  (),                                // avalon_jtag_slave.chipselect
		.av_address     (),                                //                  .address
		.av_read_n      (),                                //                  .read_n
		.av_readdata    (),                                //                  .readdata
		.av_write_n     (),                                //                  .write_n
		.av_writedata   (),                                //                  .writedata
		.av_waitrequest (),                                //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)         //               irq.irq
	);

	SEProjetoFinal_SRAM sram (
		.clk        (clk_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                  // (terminated)
	);

	SEProjetoFinal_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                          (clk_clk),                                            //                        clk_0_clk.clk
		.CPU0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                     // CPU0_reset_reset_bridge_in_reset.reset
		.CPU0_data_master_address               (cpu0_data_master_address),                           //                 CPU0_data_master.address
		.CPU0_data_master_waitrequest           (cpu0_data_master_waitrequest),                       //                                 .waitrequest
		.CPU0_data_master_byteenable            (cpu0_data_master_byteenable),                        //                                 .byteenable
		.CPU0_data_master_read                  (cpu0_data_master_read),                              //                                 .read
		.CPU0_data_master_readdata              (cpu0_data_master_readdata),                          //                                 .readdata
		.CPU0_data_master_readdatavalid         (cpu0_data_master_readdatavalid),                     //                                 .readdatavalid
		.CPU0_data_master_write                 (cpu0_data_master_write),                             //                                 .write
		.CPU0_data_master_writedata             (cpu0_data_master_writedata),                         //                                 .writedata
		.CPU0_data_master_debugaccess           (cpu0_data_master_debugaccess),                       //                                 .debugaccess
		.CPU0_instruction_master_address        (cpu0_instruction_master_address),                    //          CPU0_instruction_master.address
		.CPU0_instruction_master_waitrequest    (cpu0_instruction_master_waitrequest),                //                                 .waitrequest
		.CPU0_instruction_master_read           (cpu0_instruction_master_read),                       //                                 .read
		.CPU0_instruction_master_readdata       (cpu0_instruction_master_readdata),                   //                                 .readdata
		.CPU0_instruction_master_readdatavalid  (cpu0_instruction_master_readdatavalid),              //                                 .readdatavalid
		.CPU1_data_master_address               (cpu1_data_master_address),                           //                 CPU1_data_master.address
		.CPU1_data_master_waitrequest           (cpu1_data_master_waitrequest),                       //                                 .waitrequest
		.CPU1_data_master_byteenable            (cpu1_data_master_byteenable),                        //                                 .byteenable
		.CPU1_data_master_read                  (cpu1_data_master_read),                              //                                 .read
		.CPU1_data_master_readdata              (cpu1_data_master_readdata),                          //                                 .readdata
		.CPU1_data_master_readdatavalid         (cpu1_data_master_readdatavalid),                     //                                 .readdatavalid
		.CPU1_data_master_write                 (cpu1_data_master_write),                             //                                 .write
		.CPU1_data_master_writedata             (cpu1_data_master_writedata),                         //                                 .writedata
		.CPU1_data_master_debugaccess           (cpu1_data_master_debugaccess),                       //                                 .debugaccess
		.CPU1_instruction_master_address        (cpu1_instruction_master_address),                    //          CPU1_instruction_master.address
		.CPU1_instruction_master_waitrequest    (cpu1_instruction_master_waitrequest),                //                                 .waitrequest
		.CPU1_instruction_master_read           (cpu1_instruction_master_read),                       //                                 .read
		.CPU1_instruction_master_readdata       (cpu1_instruction_master_readdata),                   //                                 .readdata
		.CPU1_instruction_master_readdatavalid  (cpu1_instruction_master_readdatavalid),              //                                 .readdatavalid
		.CPU2_data_master_address               (cpu2_data_master_address),                           //                 CPU2_data_master.address
		.CPU2_data_master_waitrequest           (cpu2_data_master_waitrequest),                       //                                 .waitrequest
		.CPU2_data_master_byteenable            (cpu2_data_master_byteenable),                        //                                 .byteenable
		.CPU2_data_master_read                  (cpu2_data_master_read),                              //                                 .read
		.CPU2_data_master_readdata              (cpu2_data_master_readdata),                          //                                 .readdata
		.CPU2_data_master_readdatavalid         (cpu2_data_master_readdatavalid),                     //                                 .readdatavalid
		.CPU2_data_master_write                 (cpu2_data_master_write),                             //                                 .write
		.CPU2_data_master_writedata             (cpu2_data_master_writedata),                         //                                 .writedata
		.CPU2_data_master_debugaccess           (cpu2_data_master_debugaccess),                       //                                 .debugaccess
		.CPU2_instruction_master_address        (cpu2_instruction_master_address),                    //          CPU2_instruction_master.address
		.CPU2_instruction_master_waitrequest    (cpu2_instruction_master_waitrequest),                //                                 .waitrequest
		.CPU2_instruction_master_read           (cpu2_instruction_master_read),                       //                                 .read
		.CPU2_instruction_master_readdata       (cpu2_instruction_master_readdata),                   //                                 .readdata
		.CPU2_instruction_master_readdatavalid  (cpu2_instruction_master_readdatavalid),              //                                 .readdatavalid
		.CPU3_data_master_address               (cpu3_data_master_address),                           //                 CPU3_data_master.address
		.CPU3_data_master_waitrequest           (cpu3_data_master_waitrequest),                       //                                 .waitrequest
		.CPU3_data_master_byteenable            (cpu3_data_master_byteenable),                        //                                 .byteenable
		.CPU3_data_master_read                  (cpu3_data_master_read),                              //                                 .read
		.CPU3_data_master_readdata              (cpu3_data_master_readdata),                          //                                 .readdata
		.CPU3_data_master_readdatavalid         (cpu3_data_master_readdatavalid),                     //                                 .readdatavalid
		.CPU3_data_master_write                 (cpu3_data_master_write),                             //                                 .write
		.CPU3_data_master_writedata             (cpu3_data_master_writedata),                         //                                 .writedata
		.CPU3_data_master_debugaccess           (cpu3_data_master_debugaccess),                       //                                 .debugaccess
		.CPU3_instruction_master_address        (cpu3_instruction_master_address),                    //          CPU3_instruction_master.address
		.CPU3_instruction_master_waitrequest    (cpu3_instruction_master_waitrequest),                //                                 .waitrequest
		.CPU3_instruction_master_read           (cpu3_instruction_master_read),                       //                                 .read
		.CPU3_instruction_master_readdata       (cpu3_instruction_master_readdata),                   //                                 .readdata
		.CPU3_instruction_master_readdatavalid  (cpu3_instruction_master_readdatavalid),              //                                 .readdatavalid
		.CPU0_debug_mem_slave_address           (mm_interconnect_0_cpu0_debug_mem_slave_address),     //             CPU0_debug_mem_slave.address
		.CPU0_debug_mem_slave_write             (mm_interconnect_0_cpu0_debug_mem_slave_write),       //                                 .write
		.CPU0_debug_mem_slave_read              (mm_interconnect_0_cpu0_debug_mem_slave_read),        //                                 .read
		.CPU0_debug_mem_slave_readdata          (mm_interconnect_0_cpu0_debug_mem_slave_readdata),    //                                 .readdata
		.CPU0_debug_mem_slave_writedata         (mm_interconnect_0_cpu0_debug_mem_slave_writedata),   //                                 .writedata
		.CPU0_debug_mem_slave_byteenable        (mm_interconnect_0_cpu0_debug_mem_slave_byteenable),  //                                 .byteenable
		.CPU0_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu0_debug_mem_slave_waitrequest), //                                 .waitrequest
		.CPU0_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu0_debug_mem_slave_debugaccess), //                                 .debugaccess
		.CPU1_debug_mem_slave_address           (mm_interconnect_0_cpu1_debug_mem_slave_address),     //             CPU1_debug_mem_slave.address
		.CPU1_debug_mem_slave_write             (mm_interconnect_0_cpu1_debug_mem_slave_write),       //                                 .write
		.CPU1_debug_mem_slave_read              (mm_interconnect_0_cpu1_debug_mem_slave_read),        //                                 .read
		.CPU1_debug_mem_slave_readdata          (mm_interconnect_0_cpu1_debug_mem_slave_readdata),    //                                 .readdata
		.CPU1_debug_mem_slave_writedata         (mm_interconnect_0_cpu1_debug_mem_slave_writedata),   //                                 .writedata
		.CPU1_debug_mem_slave_byteenable        (mm_interconnect_0_cpu1_debug_mem_slave_byteenable),  //                                 .byteenable
		.CPU1_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu1_debug_mem_slave_waitrequest), //                                 .waitrequest
		.CPU1_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu1_debug_mem_slave_debugaccess), //                                 .debugaccess
		.CPU2_debug_mem_slave_address           (mm_interconnect_0_cpu2_debug_mem_slave_address),     //             CPU2_debug_mem_slave.address
		.CPU2_debug_mem_slave_write             (mm_interconnect_0_cpu2_debug_mem_slave_write),       //                                 .write
		.CPU2_debug_mem_slave_read              (mm_interconnect_0_cpu2_debug_mem_slave_read),        //                                 .read
		.CPU2_debug_mem_slave_readdata          (mm_interconnect_0_cpu2_debug_mem_slave_readdata),    //                                 .readdata
		.CPU2_debug_mem_slave_writedata         (mm_interconnect_0_cpu2_debug_mem_slave_writedata),   //                                 .writedata
		.CPU2_debug_mem_slave_byteenable        (mm_interconnect_0_cpu2_debug_mem_slave_byteenable),  //                                 .byteenable
		.CPU2_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu2_debug_mem_slave_waitrequest), //                                 .waitrequest
		.CPU2_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu2_debug_mem_slave_debugaccess), //                                 .debugaccess
		.CPU3_debug_mem_slave_address           (mm_interconnect_0_cpu3_debug_mem_slave_address),     //             CPU3_debug_mem_slave.address
		.CPU3_debug_mem_slave_write             (mm_interconnect_0_cpu3_debug_mem_slave_write),       //                                 .write
		.CPU3_debug_mem_slave_read              (mm_interconnect_0_cpu3_debug_mem_slave_read),        //                                 .read
		.CPU3_debug_mem_slave_readdata          (mm_interconnect_0_cpu3_debug_mem_slave_readdata),    //                                 .readdata
		.CPU3_debug_mem_slave_writedata         (mm_interconnect_0_cpu3_debug_mem_slave_writedata),   //                                 .writedata
		.CPU3_debug_mem_slave_byteenable        (mm_interconnect_0_cpu3_debug_mem_slave_byteenable),  //                                 .byteenable
		.CPU3_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu3_debug_mem_slave_waitrequest), //                                 .waitrequest
		.CPU3_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu3_debug_mem_slave_debugaccess), //                                 .debugaccess
		.SRAM_s1_address                        (mm_interconnect_0_sram_s1_address),                  //                          SRAM_s1.address
		.SRAM_s1_write                          (mm_interconnect_0_sram_s1_write),                    //                                 .write
		.SRAM_s1_readdata                       (mm_interconnect_0_sram_s1_readdata),                 //                                 .readdata
		.SRAM_s1_writedata                      (mm_interconnect_0_sram_s1_writedata),                //                                 .writedata
		.SRAM_s1_byteenable                     (mm_interconnect_0_sram_s1_byteenable),               //                                 .byteenable
		.SRAM_s1_chipselect                     (mm_interconnect_0_sram_s1_chipselect),               //                                 .chipselect
		.SRAM_s1_clken                          (mm_interconnect_0_sram_s1_clken)                     //                                 .clken
	);

	SEProjetoFinal_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu0_irq_irq)                    //    sender.irq
	);

	SEProjetoFinal_irq_mapper_001 irq_mapper_001 (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (cpu1_irq_irq)                    //    sender.irq
	);

	SEProjetoFinal_irq_mapper_001 irq_mapper_002 (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (cpu2_irq_irq)                    //    sender.irq
	);

	SEProjetoFinal_irq_mapper_001 irq_mapper_003 (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (cpu3_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (cpu0_debug_reset_request_reset),     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
