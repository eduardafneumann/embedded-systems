
module SEProjetoFinalSingle (
	clk_clk);	

	input		clk_clk;
endmodule
